module environment

@[noinit]
pub struct Environment{
	pub :
		uuid @[required] string
		
	pub 
}