module snapshot

