module environment

