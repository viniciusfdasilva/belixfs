module sys


const SYSTEM_NAME         = 'Belix'
const RELEASE_YEAR        = 2024
const AUTHOR              = 'Vinicius Silva'
const MAJOR_RELEASE       = 0
const MINOR_RELEASE       = 1

const VERSION = '${MAJOR_RELEASE.str()}.${MINOR_RELEASE.str()}' 